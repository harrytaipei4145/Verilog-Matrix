module rotation(A,rot,dir,C,clk);
input signed[35:0] A;
input dir,clk;
input [1:0] rot;

output reg signed[35:0] C;
 
//wire signed[35:0] C;
always@(posedge clk)begin
	
		if(dir==0)begin
			case(rot)
			     0:C=A;
				 1: begin C[35:32]=A[27:24];
					 C[31:28]=A[15:12];
					 C[27:24]=A[3:0];
					 C[23:20]=A[31:28];
					 C[19:16]=A[19:16];
					 C[15:12]=A[7:4];
					 C[11:8]=A[35:32];
					 C[7:4]=A[23:20];
					 C[3:0]=A[11:8];
					 end
	
				 2:	begin C[3:0]=A[35:32];
					 C[7:4]=A[31:28];
					 C[8:5]=A[27:24];
					 C[15:12]=A[23:20];
					 C[19:16]=A[19:16];
					 C[23:20]=A[15:12];
					 C[27:24]=A[11:8];
					 C[31:28]=A[7:4];
					 C[35:32]=A[3:0];
					 end
	
				 3: begin C[27:24]=A[35:32];
					 C[15:12]=A[31:28];
					 C[3:0]=A[27:24];
					 C[31:28]=A[23:20];
					 C[19:16]=A[19:16];
					 C[7:4]=A[15:12];
					 C[35:32]=A[11:8];
					 C[23:20]=A[7:4];
					 C[11:8]=A[3:0];
					 end
	
			endcase	 
		end


		else begin
			case(rot)
			0:C=A;
				 1: begin C[27:24]=A[35:32];
					 C[15:12]=A[31:28];
					 C[3:0]=A[27:24];
					 C[31:28]=A[23:20];
					 C[19:16]=A[19:16];
					 C[7:4]=A[15:12];
					 C[35:32]=A[11:8];
					 C[23:20]=A[7:4];
					 C[11:8]=A[3:0];
					 end
	
				2:begin   C[35:32]=A[3:0];
					 C[31:28]=A[7:4];
					 C[27:24]=A[8:5];
					 C[23:20]=A[15:12];
					 C[19:16]=A[19:16];
					 C[15:12]=A[23:20];
					 C[11:8]=A[27:24];
					 C[7:4]=A[31:28];
					 C[3:0]=A[35:32];
				end
	
				3:begin   C[35:32]=A[27:24];
					 C[31:28]=A[15:12];
					 C[27:24]=A[3:0];
					 C[23:20]=A[31:28];
					 C[19:16]=A[19:16];
					 C[15:12]=A[7:4];
					 C[11:8]=A[35:32];
					 C[7:4]=A[23:20];
					 C[3:0]=A[11:8];
					 end
	
			endcase
		end
	
end
endmodule